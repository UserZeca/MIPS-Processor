library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all; -- Corrigido (removido std_logic_arith)

entity LZCShifter_28_to_28_counting_32_comb_uid16 is
    port ( I : in  std_logic_vector(27 downto 0);
           Count : out  std_logic_vector(4 downto 0);
           O : out  std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_comb_uid16 is
signal level5 :  std_logic_vector(27 downto 0);
signal count4 :  std_logic;
signal level4 :  std_logic_vector(27 downto 0);
signal count3 :  std_logic;
signal level3 :  std_logic_vector(27 downto 0);
signal count2 :  std_logic;
signal level2 :  std_logic_vector(27 downto 0);
signal count1 :  std_logic;
signal level1 :  std_logic_vector(27 downto 0);
signal count0 :  std_logic;
signal level0 :  std_logic_vector(27 downto 0);
signal sCount :  std_logic_vector(4 downto 0);
begin
    level5 <= I ;
    count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
    level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

    count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
    level3<= level4(27 downto 0) when count3='0' else level4(19 downto 0) & (7 downto 0 => '0');

    count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
    level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

    count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
    level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

    count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
    level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

    O <= level0;
    sCount <= count4 & count3 & count2 & count1 & count0;
    Count <= sCount;
end architecture;